module floatadd #(
    parameters
) (
    input [15:0] a, // 16-bit floating point input a
    input [15:0] b, // 16-bit floating point input b
    output [15:0] result // 16-bit floating point output result
);

reg sign;
reg 


endmodule