module convolve (
    ports
);
    
endmodule